Library IEEE;
	use IEEE.std_logic_1164.all;
entity testing is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A43: buffer std_logic
);
end testing;

architecture testing_behav of testing is
signal n_32,n_33,n_37,n_38,n_39,n_40,n_46,n_47,n_48,n_49,n_55,n_56,n_57,n_58,n_59,n_60,n_66,n_67,n_68,n_69,n_72,n_73,n_74,n_81,n_82,n_83,n_84,n_87,n_88,n_91,n_94,n_97,n_98,n_99,n_104,n_105,n_106,n_107,n_108,n_109,n_114,n_120,n_121,n_122,n_123,n_126,n_127,n_128,n_129,n_130,n_135,n_136,n_140,n_141,n_142,n_143,n_149,n_150,n_151,n_152,n_158,n_159,n_160,n_161,n_166,n_167,n_171,n_172,n_173,n_174,n_180,n_181,n_182,n_183,n_189,n_190,n_191,n_192,n_193,n_194,n_195,n_196,n_197,n_201,n_204,n_207,n_208,n_209,n_214,n_215,n_216,n_217,n_218,n_223,n_224,n_225,n_226,n_227,n_234,n_235,n_239,n_240,n_241,n_242,n_248,n_249,n_250,n_251,n_257,n_258,n_259,n_260,n_261,n_262,n_265,n_268,n_271,n_272,n_275,n_278,n_281,n_282,n_283,n_288,n_289,n_290,n_291,n_292,n_293,n_298,n_301,n_304,n_307,n_308,n_309,n_314,n_315,n_316,n_317,n_318,n_319,n_320,n_321,n_322,n_323,n_328,n_333,n_334,n_338,n_339,n_340,n_341,n_347,n_348,n_349,n_350,n_356,n_357,n_358,n_359,n_360,n_361,n_364,n_367,n_370,n_371,n_372,n_377,n_378,n_379,n_380,n_381,n_382,n_383,n_384,n_385,n_386,n_391,n_397,n_398,n_402,n_403,n_404,n_405,n_411,n_412,n_413,n_414,n_420,n_421,n_422,n_423,n_424,n_425,n_428,n_431,n_434,n_435,n_436,n_441,n_442,n_443,n_444,n_445,n_446,n_451,n_456,n_457,n_461,n_462,n_463,n_464,n_470,n_471,n_472,n_473,n_479,n_480,n_481,n_482,n_483,n_484,n_485,n_486,n_487,n_488,n_489,n_490,n_491,n_492,n_493,n_494,n_495,n_496: std_logic;
begin

A43 <=( (not n_496) );
 n_32 <=( (not A202)  and  A203 );
 n_33 <=( A200  and  n_32 );
 n_37 <=( A202  and  (not A203) );
 n_38 <=( (not A200)  and  n_37 );
 n_39 <=( n_38 ) or ( n_33 );
 n_40 <=( (not A199)  and  n_39 );
 n_46 <=( A202  and  (not A203) );
 n_47 <=( A199  and  n_46 );
 n_48 <=( n_47 ) or ( A201 );
 n_49 <=( A200  and  n_48 );
 n_55 <=( (not A202)  and  A203 );
 n_56 <=( (not A200)  and  n_55 );
 n_57 <=( n_56 ) or ( A201 );
 n_58 <=( A199  and  n_57 );
 n_59 <=( n_58 ) or ( n_49 );
 n_60 <=( n_59 ) or ( n_40 );
 n_66 <=( A170 ) or ( A169 );
 n_67 <=( A168  and  n_66 );
 n_68 <=( (not A167)  and  n_67 );
 n_69 <=( A166  and  n_68 );
 n_72 <=( (not A166)  and  A167 );
 n_73 <=( n_72 ) or ( n_69 );
 n_74 <=( n_60  and  n_73 );
 n_81 <=( (not A169)  and  (not A170) );
 n_82 <=( n_81 ) or ( (not A168) );
 n_83 <=( n_82 ) or ( (not A166) );
 n_84 <=( (not A167)  and  n_83 );
 n_87 <=( A166  and  A167 );
 n_88 <=( n_87 ) or ( n_84 );
 n_91 <=( (not A203) ) or ( A202 );
 n_94 <=( (not A199)  and  A200 );
 n_97 <=( A199  and  (not A200) );
 n_98 <=( n_97 ) or ( n_94 );
 n_99 <=( n_91  and  n_98 );
 n_104 <=( A203 ) or ( (not A202) );
 n_105 <=( A200  and  n_104 );
 n_106 <=( A199  and  n_105 );
 n_107 <=( n_106 ) or ( n_99 );
 n_108 <=( n_88  and  n_107 );
 n_109 <=( (not A201)  and  n_108 );
 n_114 <=( A203 ) or ( (not A202) );
 n_120 <=( (not A169)  and  (not A170) );
 n_121 <=( n_120 ) or ( (not A168) );
 n_122 <=( n_121 ) or ( (not A166) );
 n_123 <=( (not A167)  and  n_122 );
 n_126 <=( A166  and  A167 );
 n_127 <=( n_126 ) or ( n_123 );
 n_128 <=( n_114  and  n_127 );
 n_129 <=( (not A200)  and  n_128 );
 n_130 <=( (not A199)  and  n_129 );
 n_135 <=( (not A268)  and  A269 );
 n_136 <=( A266  and  n_135 );
 n_140 <=( A268  and  (not A269) );
 n_141 <=( (not A266)  and  n_140 );
 n_142 <=( n_141 ) or ( n_136 );
 n_143 <=( (not A265)  and  n_142 );
 n_149 <=( A268  and  (not A269) );
 n_150 <=( A265  and  n_149 );
 n_151 <=( n_150 ) or ( A267 );
 n_152 <=( A266  and  n_151 );
 n_158 <=( (not A268)  and  A269 );
 n_159 <=( (not A266)  and  n_158 );
 n_160 <=( n_159 ) or ( A267 );
 n_161 <=( A265  and  n_160 );
 n_166 <=( (not A301)  and  A302 );
 n_167 <=( A299  and  n_166 );
 n_171 <=( A301  and  (not A302) );
 n_172 <=( (not A299)  and  n_171 );
 n_173 <=( n_172 ) or ( n_167 );
 n_174 <=( (not A298)  and  n_173 );
 n_180 <=( A301  and  (not A302) );
 n_181 <=( A298  and  n_180 );
 n_182 <=( n_181 ) or ( A300 );
 n_183 <=( A299  and  n_182 );
 n_189 <=( (not A301)  and  A302 );
 n_190 <=( (not A299)  and  n_189 );
 n_191 <=( n_190 ) or ( A300 );
 n_192 <=( A298  and  n_191 );
 n_193 <=( n_192 ) or ( n_183 );
 n_194 <=( n_193 ) or ( n_174 );
 n_195 <=( n_194 ) or ( n_161 );
 n_196 <=( n_195 ) or ( n_152 );
 n_197 <=( n_196 ) or ( n_143 );
 n_201 <=( (not A236) ) or ( A235 );
 n_204 <=( (not A232)  and  A233 );
 n_207 <=( A232  and  (not A233) );
 n_208 <=( n_207 ) or ( n_204 );
 n_209 <=( n_201  and  n_208 );
 n_214 <=( A236 ) or ( (not A235) );
 n_215 <=( A233  and  n_214 );
 n_216 <=( A232  and  n_215 );
 n_217 <=( n_216 ) or ( n_209 );
 n_218 <=( (not A234)  and  n_217 );
 n_223 <=( A236 ) or ( (not A235) );
 n_224 <=( (not A233)  and  n_223 );
 n_225 <=( (not A232)  and  n_224 );
 n_226 <=( n_225 ) or ( n_218 );
 n_227 <=( n_197  and  n_226 );
 n_234 <=( (not A235)  and  A236 );
 n_235 <=( A233  and  n_234 );
 n_239 <=( A235  and  (not A236) );
 n_240 <=( (not A233)  and  n_239 );
 n_241 <=( n_240 ) or ( n_235 );
 n_242 <=( (not A232)  and  n_241 );
 n_248 <=( A235  and  (not A236) );
 n_249 <=( A232  and  n_248 );
 n_250 <=( n_249 ) or ( A234 );
 n_251 <=( A233  and  n_250 );
 n_257 <=( (not A235)  and  A236 );
 n_258 <=( (not A233)  and  n_257 );
 n_259 <=( n_258 ) or ( A234 );
 n_260 <=( A232  and  n_259 );
 n_261 <=( n_260 ) or ( n_251 );
 n_262 <=( n_261 ) or ( n_242 );
 n_265 <=( (not A302) ) or ( A301 );
 n_268 <=( (not A298)  and  A299 );
 n_271 <=( A298  and  (not A299) );
 n_272 <=( n_271 ) or ( n_268 );
 n_275 <=( (not A269) ) or ( A268 );
 n_278 <=( (not A265)  and  A266 );
 n_281 <=( A265  and  (not A266) );
 n_282 <=( n_281 ) or ( n_278 );
 n_283 <=( n_275  and  n_282 );
 n_288 <=( A269 ) or ( (not A268) );
 n_289 <=( A266  and  n_288 );
 n_290 <=( A265  and  n_289 );
 n_291 <=( n_290 ) or ( n_283 );
 n_292 <=( n_272  and  n_291 );
 n_293 <=( n_265  and  n_292 );
 n_298 <=( A302 ) or ( (not A301) );
 n_301 <=( (not A269) ) or ( A268 );
 n_304 <=( (not A265)  and  A266 );
 n_307 <=( A265  and  (not A266) );
 n_308 <=( n_307 ) or ( n_304 );
 n_309 <=( n_301  and  n_308 );
 n_314 <=( A269 ) or ( (not A268) );
 n_315 <=( A266  and  n_314 );
 n_316 <=( A265  and  n_315 );
 n_317 <=( n_316 ) or ( n_309 );
 n_318 <=( n_298  and  n_317 );
 n_319 <=( A299  and  n_318 );
 n_320 <=( A298  and  n_319 );
 n_321 <=( n_320 ) or ( n_293 );
 n_322 <=( n_262  and  n_321 );
 n_323 <=( (not A267)  and  n_322 );
 n_328 <=( A269 ) or ( (not A268) );
 n_333 <=( (not A235)  and  A236 );
 n_334 <=( A233  and  n_333 );
 n_338 <=( A235  and  (not A236) );
 n_339 <=( (not A233)  and  n_338 );
 n_340 <=( n_339 ) or ( n_334 );
 n_341 <=( (not A232)  and  n_340 );
 n_347 <=( A235  and  (not A236) );
 n_348 <=( A232  and  n_347 );
 n_349 <=( n_348 ) or ( A234 );
 n_350 <=( A233  and  n_349 );
 n_356 <=( (not A235)  and  A236 );
 n_357 <=( (not A233)  and  n_356 );
 n_358 <=( n_357 ) or ( A234 );
 n_359 <=( A232  and  n_358 );
 n_360 <=( n_359 ) or ( n_350 );
 n_361 <=( n_360 ) or ( n_341 );
 n_364 <=( (not A302) ) or ( A301 );
 n_367 <=( (not A298)  and  A299 );
 n_370 <=( A298  and  (not A299) );
 n_371 <=( n_370 ) or ( n_367 );
 n_372 <=( n_364  and  n_371 );
 n_377 <=( A302 ) or ( (not A301) );
 n_378 <=( A299  and  n_377 );
 n_379 <=( A298  and  n_378 );
 n_380 <=( n_379 ) or ( n_372 );
 n_381 <=( n_361  and  n_380 );
 n_382 <=( n_328  and  n_381 );
 n_383 <=( (not A266)  and  n_382 );
 n_384 <=( (not A265)  and  n_383 );
 n_385 <=( n_384 ) or ( n_323 );
 n_386 <=( (not A300)  and  n_385 );
 n_391 <=( A302 ) or ( (not A301) );
 n_397 <=( (not A235)  and  A236 );
 n_398 <=( A233  and  n_397 );
 n_402 <=( A235  and  (not A236) );
 n_403 <=( (not A233)  and  n_402 );
 n_404 <=( n_403 ) or ( n_398 );
 n_405 <=( (not A232)  and  n_404 );
 n_411 <=( A235  and  (not A236) );
 n_412 <=( A232  and  n_411 );
 n_413 <=( n_412 ) or ( A234 );
 n_414 <=( A233  and  n_413 );
 n_420 <=( (not A235)  and  A236 );
 n_421 <=( (not A233)  and  n_420 );
 n_422 <=( n_421 ) or ( A234 );
 n_423 <=( A232  and  n_422 );
 n_424 <=( n_423 ) or ( n_414 );
 n_425 <=( n_424 ) or ( n_405 );
 n_428 <=( (not A269) ) or ( A268 );
 n_431 <=( (not A265)  and  A266 );
 n_434 <=( A265  and  (not A266) );
 n_435 <=( n_434 ) or ( n_431 );
 n_436 <=( n_428  and  n_435 );
 n_441 <=( A269 ) or ( (not A268) );
 n_442 <=( A266  and  n_441 );
 n_443 <=( A265  and  n_442 );
 n_444 <=( n_443 ) or ( n_436 );
 n_445 <=( n_425  and  n_444 );
 n_446 <=( (not A267)  and  n_445 );
 n_451 <=( A269 ) or ( (not A268) );
 n_456 <=( (not A235)  and  A236 );
 n_457 <=( A233  and  n_456 );
 n_461 <=( A235  and  (not A236) );
 n_462 <=( (not A233)  and  n_461 );
 n_463 <=( n_462 ) or ( n_457 );
 n_464 <=( (not A232)  and  n_463 );
 n_470 <=( A235  and  (not A236) );
 n_471 <=( A232  and  n_470 );
 n_472 <=( n_471 ) or ( A234 );
 n_473 <=( A233  and  n_472 );
 n_479 <=( (not A235)  and  A236 );
 n_480 <=( (not A233)  and  n_479 );
 n_481 <=( n_480 ) or ( A234 );
 n_482 <=( A232  and  n_481 );
 n_483 <=( n_482 ) or ( n_473 );
 n_484 <=( n_483 ) or ( n_464 );
 n_485 <=( n_451  and  n_484 );
 n_486 <=( (not A266)  and  n_485 );
 n_487 <=( (not A265)  and  n_486 );
 n_488 <=( n_487 ) or ( n_446 );
 n_489 <=( n_391  and  n_488 );
 n_490 <=( (not A299)  and  n_489 );
 n_491 <=( (not A298)  and  n_490 );
 n_492 <=( n_491 ) or ( n_386 );
 n_493 <=( n_492 ) or ( n_227 );
 n_494 <=( n_493 ) or ( n_130 );
 n_495 <=( n_494 ) or ( n_109 );
 n_496 <=( n_495 ) or ( n_74 );


end testing_behav;
