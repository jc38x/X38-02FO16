Library IEEE;
	use IEEE.std_logic_1164.all;
entity testing is
	Port (
	A302,A301,A300,A299,A298,A269,A268,A267,A266,A265,A236,A235,A234,A233,A232,A203,A202,A201,A200,A199,A166,A167,A168,A169,A170: in std_logic;
	A142,A141,A140,A139,A138,A109,A108,A107,A106,A105,A76,A75,A74,A73,A72,A43,A42,A41,A40,A39,A6,A7,A8,A9,A10: buffer std_logic
);
end testing;

architecture testing_behav of testing is
signal a50a,a51a,a52a,a53a,a54a,a55a,a56a,a57a,a58a,a59a,a60a,a61a,a62a,a63a,a64a,a65a,a66a,a67a,a68a,a69a,a70a,a71a,a72a,a73a,a74a,a75a,a76a,a77a,a78a,a79a,a80a,a81a,a82a,a83a,a84a,a85a,a86a,a87a,a88a,a89a,a90a,a91a,a92a,a93a,a94a,a95a,a96a,a97a,a98a,a99a,a100a,a101a,a102a,a103a,a104a,a105a,a106a,a107a,a108a,a109a,a110a,a111a,a112a,a113a,a114a,a115a,a116a,a117a,a118a,a119a,a120a,a121a,a122a,a123a,a124a,a125a,a126a,a127a,a128a,a129a,a130a,a131a,a132a,a133a,a134a,a135a,a136a,a137a,a138a,a139a,a140a,a141a,a142a,a143a,a144a,a145a,a146a,a147a,a148a,a149a,a150a,a151a,a152a,a153a,a154a,a155a,a156a,a157a,a158a,a160a,a161a,a162a,a163a,a164a,a165a,a166a,a167a,a168a,a169a,a170a,a171a,a173a,a174a,a175a,a176a,a177a,a178a,a179a,a180a,a181a,a182a,a183a,a184a,a185a,a186a,a187a,a188a,a189a,a190a,a191a,a192a,a193a,a194a,a195a,a196a,a197a,a198a,a199a,a200a,a201a,a202a,a203a,a204a,a205a,a206a,a207a,a208a,a209a,a210a,a211a,a212a,a213a,a214a,a215a,a216a,a217a,a218a,a219a,a220a,a221a,a222a,a223a,a224a,a225a,a226a,a227a,a228a,a229a,a230a,a231a,a232a,a233a,a234a,a235a,a236a,a237a,a238a,a239a,a240a,a241a,a242a,a243a,a244a,a245a,a246a,a247a,a248a,a249a,a250a,a252a,a253a,a254a,a255a,a256a,a257a,a258a,a259a,a260a,a261a,a262a,a263a,a264a,a265a,a266a,a267a,a268a,a269a,a270a,a271a,a272a,a273a,a274a,a275a,a276a,a277a,a278a,a279a,a280a,a281a,a282a,a283a,a284a,a285a,a286a,a287a,a288a,a289a,a290a,a291a,a292a,a293a,a294a,a295a,a296a,a297a,a298a,a299a,a300a,a301a,a302a,a303a,a304a,a305a,a306a,a307a,a308a,a309a,a310a,a311a,a312a,a314a,a315a,a316a,a317a,a318a,a320a,a321a,a322a,a323a,a324a,a325a,a326a,a327a,a328a,a329a,a330a,a331a,a332a,a333a,a334a,a335a,a336a,a337a,a338a,a339a,a340a,a341a,a342a,a343a,a344a,a345a,a346a,a347a,a348a,a349a,a350a,a351a,a352a,a354a,a355a,a356a,a357a,a358a,a359a,a360a,a361a,a362a,a363a,a364a,a365a,a366a,a367a,a368a,a369a,a370a,a371a,a372a,a373a,a374a,a375a,a376a,a377a,a378a,a379a,a380a,a381a,a382a,a383a,a384a,a385a,a386a,a387a,a388a,a389a,a390a,a391a,a392a,a393a,a394a,a395a,a396a,a397a,a398a,a399a,a400a,a401a,a402a,a403a,a404a,a406a,a407a,a408a,a409a,a410a,a412a,a413a,a414a,a415a,a416a,a417a,a418a,a419a,a420a,a421a,a422a,a423a,a424a,a425a,a426a,a427a,a428a,a429a,a430a,a431a,a432a,a433a,a434a,a435a,a436a,a437a,a438a,a439a,a440a,a441a,a442a,a443a,a444a,a445a,a446a,a447a,a448a,a449a,a450a,a451a,a452a,a453a,a454a,a455a,a457a,a458a,a459a,a460a,a461a,a462a,a463a,a464a,a465a,a466a,a467a,a468a,a469a,a470a,a471a,a472a,a473a,a474a,a475a,a476a,a477a,a478a,a479a,a480a,a481a,a482a,a483a,a484a,a485a,a486a,a487a,a488a,a489a,a490a,a491a,a492a,a493a,a494a,a495a,a496a,a497a,a498a,a499a,a500a,a501a,a502a,a503a,a504a,a505a,a506a,a507a,a508a,a509a,a510a,a511a,a512a,a513a,a514a,a515a,a516a,a517a,a518a,a519a,a520a,a521a,a522a,a523a,a524a,a525a,a526a,a527a,a528a,a529a,a530a,a531a,a532a,a533a,a534a,a535a,a536a,a538a,a539a,a540a,a541a,a542a,a543a,a544a,a545a,a546a,a547a,a548a,a549a,a550a,a552a,a553a,a554a,a555a,a556a,a557a,a558a,a559a,a560a,a561a,a562a,a563a,a564a,a565a,a566a,a567a,a568a,a569a,a570a,a571a,a572a,a573a,a574a,a575a,a576a,a577a,a578a,a579a,a580a,a581a,a582a,a583a,a584a,a585a,a586a,a587a,a588a,a589a,a590a,a591a,a592a,a593a,a594a,a595a,a596a,a597a,a598a,a599a,a600a,a601a,a602a,a603a,a604a,a605a,a606a,a607a,a608a,a609a,a610a,a611a,a612a,a613a,a614a,a615a,a616a,a617a,a618a,a619a,a620a,a621a,a622a,a623a,a624a,a625a,a626a,a627a,a628a,a629a,a630a,a631a,a632a,a633a,a634a,a635a,a636a,a637a,a638a,a639a,a640a,a641a,a642a,a643a,a644a,a645a,a646a,a647a,a648a,a649a,a650a,a651a,a652a,a653a,a654a,a656a,a657a,a658a,a659a,a660a,a661a,a662a,a663a,a664a,a665a,a666a,a667a,a668a,a669a,a670a,a671a,a672a,a673a,a674a,a675a,a676a,a677a,a678a,a679a,a680a,a681a,a682a,a683a,a684a,a685a,a686a,a687a,a688a,a689a,a690a,a691a,a692a,a693a,a694a,a695a,a696a,a697a,a698a,a699a,a700a,a701a,a702a,a703a,a704a,a705a,a706a,a707a,a708a,a709a,a710a,a711a,a712a,a713a,a714a,a715a,a716a,a717a,a718a,a719a,a720a,a721a,a722a,a723a,a724a,a725a,a726a,a727a,a728a,a729a,a730a,a731a,a732a,a733a,a734a,a736a,a737a,a738a,a739a,a740a,a741a,a742a,a743a,a744a,a745a,a746a,a747a,a748a,a749a,a750a,a751a,a752a,a753a,a754a,a755a,a756a,a757a,a758a,a759a,a760a,a761a,a762a,a763a,a764a,a765a,a766a,a767a,a768a,a769a,a770a,a771a,a772a,a773a,a774a,a775a,a776a,a777a,a778a,a779a,a780a,a781a,a782a,a783a,a784a,a785a,a786a,a787a,a788a,a789a,a790a,a791a,a792a,a793a,a794a,a795a,a796a,a797a,a798a,a799a,a800a,a801a,a802a,a803a,a804a,a805a,a806a,a808a,a809a,a810a,a811a,a812a,a813a,a814a,a815a,a816a,a817a,a818a,a819a,a820a,a821a,a822a,a823a,a824a,a825a,a826a,a827a,a828a,a829a,a830a,a831a,a832a,a833a,a834a,a835a,a836a,a837a,a839a,a840a,a841a,a842a,a843a,a844a,a845a,a846a,a847a,a848a,a849a,a850a,a851a,a852a,a853a: std_logic;
begin

a50a <=( (not A169)  and  A170 );
 a51a <=( (not A166)  and  A167 );
 a52a <=( A166  and  (not A167) );
 a53a <=( (not a51a)  and  (not a52a) );
 a54a <=( (not A200)  and  A199 );
 a55a <=( A200  and  (not A199) );
 a56a <=( (not a54a)  and  (not a55a) );
 a57a <=( (not A203)  and  (not A202) );
 a58a <=( A201  and  (not a57a) );
 a59a <=( (not A203)  and  (not A201) );
 a60a <=( (not A202)  and  a59a );
 a61a <=( (not a58a)  and  (not a60a) );
 a62a <=( (not a56a)  and  (not a61a) );
 a63a <=( A168  and  (not a53a) );
 a64a <=( a62a  and  a63a );
 a65a <=( (not A201)  and  (not a57a) );
 a66a <=( (not A203)  and  A201 );
 a67a <=( (not A202)  and  a66a );
 a68a <=( A200  and  A199 );
 a69a <=( (not A200)  and  (not A199) );
 a70a <=( (not a68a)  and  (not a69a) );
 a71a <=( (not a67a)  and  a70a );
 a72a <=( (not a65a)  and  a71a );
 a73a <=( (not A168)  and  (not a72a) );
 a74a <=( (not a64a)  and  (not a73a) );
 a75a <=( (not a50a)  and  (not a74a) );
 a76a <=( (not a53a)  and  (not a56a) );
 a77a <=( A201  and  (not A168) );
 a78a <=( a76a  and  a77a );
 a79a <=( (not A201)  and  A168 );
 a80a <=( (not a78a)  and  (not a79a) );
 a81a <=( a50a  and  (not a80a) );
 a82a <=( A166  and  A167 );
 a83a <=( (not A166)  and  (not A167) );
 a84a <=( (not a82a)  and  (not a83a) );
 a85a <=( (not A201)  and  (not a84a) );
 a86a <=( (not a81a)  and  (not a85a) );
 a87a <=( (not a57a)  and  (not a86a) );
 a88a <=( A168  and  a50a );
 a89a <=( a84a  and  (not a88a) );
 a90a <=( (not a71a)  and  (not a89a) );
 a91a <=( (not A201)  and  (not A168) );
 a92a <=( a57a  and  a91a );
 a93a <=( a50a  and  a92a );
 a94a <=( a76a  and  a93a );
 a95a <=( (not A236)  and  (not A235) );
 a96a <=( A299  and  (not A298) );
 a97a <=( (not A299)  and  A298 );
 a98a <=( (not a96a)  and  (not a97a) );
 a99a <=( (not A302)  and  (not A301) );
 a100a <=( A300  and  (not a99a) );
 a101a <=( (not A302)  and  (not A300) );
 a102a <=( (not A301)  and  a101a );
 a103a <=( (not a100a)  and  (not a102a) );
 a104a <=( (not a98a)  and  (not a103a) );
 a105a <=( A266  and  (not A265) );
 a106a <=( (not A266)  and  A265 );
 a107a <=( (not a105a)  and  (not a106a) );
 a108a <=( (not A269)  and  (not A268) );
 a109a <=( A267  and  (not a108a) );
 a110a <=( (not A269)  and  (not A267) );
 a111a <=( (not A268)  and  a110a );
 a112a <=( (not a109a)  and  (not a111a) );
 a113a <=( (not a107a)  and  (not a112a) );
 a114a <=( (not a104a)  and  (not a113a) );
 a115a <=( (not A234)  and  (not a114a) );
 a116a <=( (not A233)  and  A232 );
 a117a <=( A233  and  (not A232) );
 a118a <=( (not a116a)  and  (not a117a) );
 a119a <=( (not A267)  and  (not a108a) );
 a120a <=( (not A269)  and  A267 );
 a121a <=( (not A268)  and  a120a );
 a122a <=( A266  and  A265 );
 a123a <=( (not A266)  and  (not A265) );
 a124a <=( (not a122a)  and  (not a123a) );
 a125a <=( (not a121a)  and  a124a );
 a126a <=( (not a119a)  and  a125a );
 a127a <=( (not A300)  and  (not a99a) );
 a128a <=( (not A302)  and  A300 );
 a129a <=( (not A301)  and  a128a );
 a130a <=( A299  and  A298 );
 a131a <=( (not A299)  and  (not A298) );
 a132a <=( (not a130a)  and  (not a131a) );
 a133a <=( (not a129a)  and  a132a );
 a134a <=( (not a127a)  and  a133a );
 a135a <=( (not a126a)  and  (not a134a) );
 a136a <=( (not a118a)  and  a135a );
 a137a <=( A234  and  a136a );
 a138a <=( (not a115a)  and  (not a137a) );
 a139a <=( (not a95a)  and  (not a138a) );
 a140a <=( (not A236)  and  A234 );
 a141a <=( (not A235)  and  a140a );
 a142a <=( A233  and  A232 );
 a143a <=( (not A233)  and  (not A232) );
 a144a <=( (not a142a)  and  (not a143a) );
 a145a <=( (not a141a)  and  a144a );
 a146a <=( (not a98a)  and  (not a145a) );
 a147a <=( (not a103a)  and  a146a );
 a148a <=( (not a107a)  and  (not a145a) );
 a149a <=( (not a112a)  and  a148a );
 a150a <=( (not A236)  and  (not A234) );
 a151a <=( (not A235)  and  a150a );
 a152a <=( a136a  and  a151a );
 a153a <=( (not a90a)  and  (not a94a) );
 a154a <=( (not a149a)  and  a153a );
 a155a <=( (not a147a)  and  a154a );
 a156a <=( (not a152a)  and  a155a );
 a157a <=( (not a75a)  and  a156a );
 a158a <=( (not a87a)  and  a157a );
 A142 <=( (not a139a)  and  a158a );
 a160a <=( A168  and  (not a50a) );
 a161a <=( (not A168)  and  a50a );
 a162a <=( (not a160a)  and  (not a161a) );
 a163a <=( (not A234)  and  (not a95a) );
 a164a <=( a145a  and  (not a163a) );
 a165a <=( (not a62a)  and  a164a );
 a166a <=( (not a135a)  and  a165a );
 a167a <=( (not a53a)  and  (not a162a) );
 a168a <=( (not a166a)  and  a167a );
 a169a <=( (not A168)  and  (not a50a) );
 a170a <=( a89a  and  (not a169a) );
 a171a <=( (not a72a)  and  (not a170a) );
 A141 <=( (not a168a)  and  (not a171a) );
 a173a <=( A234  and  (not a95a) );
 a174a <=( (not a151a)  and  (not a173a) );
 a175a <=( (not a118a)  and  (not a174a) );
 a176a <=( (not a61a)  and  a175a );
 a177a <=( (not a61a)  and  a104a );
 a178a <=( (not a170a)  and  a177a );
 a179a <=( (not a176a)  and  (not a178a) );
 a180a <=( (not a56a)  and  (not a179a) );
 a181a <=( (not a162a)  and  a175a );
 a182a <=( a104a  and  (not a162a) );
 a183a <=( (not a72a)  and  a182a );
 a184a <=( (not a181a)  and  (not a183a) );
 a185a <=( (not a53a)  and  (not a184a) );
 a186a <=( (not a113a)  and  (not a185a) );
 a187a <=( (not a180a)  and  a186a );
 a188a <=( (not A267)  and  (not A168) );
 a189a <=( a104a  and  a188a );
 a190a <=( A168  and  (not a107a) );
 a191a <=( (not a53a)  and  a190a );
 a192a <=( (not a134a)  and  a191a );
 a193a <=( A267  and  a192a );
 a194a <=( (not a189a)  and  (not a193a) );
 a195a <=( (not a108a)  and  (not a194a) );
 a196a <=( (not A168)  and  (not a98a) );
 a197a <=( (not a125a)  and  a196a );
 a198a <=( (not a103a)  and  a197a );
 a199a <=( a111a  and  a192a );
 a200a <=( (not a198a)  and  (not a199a) );
 a201a <=( (not a195a)  and  a200a );
 a202a <=( (not a50a)  and  (not a201a) );
 a203a <=( (not a89a)  and  a104a );
 a204a <=( (not a126a)  and  a203a );
 a205a <=( (not a107a)  and  a161a );
 a206a <=( (not a53a)  and  a205a );
 a207a <=( (not a112a)  and  a206a );
 a208a <=( (not a134a)  and  a207a );
 a209a <=( (not a204a)  and  (not a208a) );
 a210a <=( (not a202a)  and  a209a );
 a211a <=( (not a61a)  and  (not a210a) );
 a212a <=( (not a176a)  and  (not a211a) );
 a213a <=( (not a56a)  and  (not a212a) );
 a214a <=( (not a72a)  and  (not a126a) );
 a215a <=( a182a  and  a214a );
 a216a <=( (not a181a)  and  (not a215a) );
 a217a <=( (not a53a)  and  (not a216a) );
 a218a <=( a113a  and  (not a134a) );
 a219a <=( a171a  and  a218a );
 a220a <=( (not a217a)  and  (not a219a) );
 a221a <=( (not a213a)  and  a220a );
 a222a <=( (not a98a)  and  (not a118a) );
 a223a <=( (not a126a)  and  a222a );
 a224a <=( A234  and  a223a );
 a225a <=( A300  and  a224a );
 a226a <=( (not A300)  and  (not A234) );
 a227a <=( (not a225a)  and  (not a226a) );
 a228a <=( (not a99a)  and  (not a227a) );
 a229a <=( (not A300)  and  a224a );
 a230a <=( A300  and  (not A234) );
 a231a <=( (not a229a)  and  (not a230a) );
 a232a <=( a99a  and  (not a231a) );
 a233a <=( (not a113a)  and  a132a );
 a234a <=( (not A234)  and  (not a233a) );
 a235a <=( (not a232a)  and  (not a234a) );
 a236a <=( (not a228a)  and  a235a );
 a237a <=( (not a95a)  and  (not a236a) );
 a238a <=( (not A300)  and  (not a145a) );
 a239a <=( a151a  and  a223a );
 a240a <=( A300  and  a239a );
 a241a <=( (not a238a)  and  (not a240a) );
 a242a <=( (not a99a)  and  (not a241a) );
 a243a <=( (not a113a)  and  a133a );
 a244a <=( (not a145a)  and  (not a243a) );
 a245a <=( a102a  and  a239a );
 a246a <=( a153a  and  (not a244a) );
 a247a <=( (not a245a)  and  a246a );
 a248a <=( (not a75a)  and  a247a );
 a249a <=( (not a87a)  and  a248a );
 a250a <=( (not a242a)  and  a249a );
 A138 <=( (not a237a)  and  a250a );
 a252a <=( A234  and  (not A233) );
 a253a <=( (not a95a)  and  a252a );
 a254a <=( A232  and  (not a253a) );
 a255a <=( (not a143a)  and  (not a254a) );
 a256a <=( A300  and  a97a );
 a257a <=( (not a99a)  and  a256a );
 a258a <=( A267  and  a106a );
 a259a <=( (not a108a)  and  a258a );
 a260a <=( (not a96a)  and  (not a105a) );
 a261a <=( (not a259a)  and  a260a );
 a262a <=( (not a257a)  and  a261a );
 a263a <=( (not a255a)  and  (not a262a) );
 a264a <=( A169  and  (not A170) );
 a265a <=( (not A167)  and  a264a );
 a266a <=( A167  and  a50a );
 a267a <=( (not a265a)  and  (not a266a) );
 a268a <=( (not A166)  and  (not a267a) );
 a269a <=( A166  and  a264a );
 a270a <=( (not A168)  and  (not a269a) );
 a271a <=( A167  and  (not a270a) );
 a272a <=( (not A167)  and  a50a );
 a273a <=( (not A168)  and  (not a272a) );
 a274a <=( A166  and  (not a273a) );
 a275a <=( (not a271a)  and  (not a274a) );
 a276a <=( (not a268a)  and  a275a );
 a277a <=( A201  and  a54a );
 a278a <=( (not a57a)  and  a277a );
 a279a <=( (not a55a)  and  (not a278a) );
 a280a <=( (not a276a)  and  (not a279a) );
 a281a <=( A201  and  (not A200) );
 a282a <=( (not a57a)  and  a281a );
 a283a <=( A199  and  (not a282a) );
 a284a <=( (not a69a)  and  (not a283a) );
 a285a <=( (not A167)  and  A169 );
 a286a <=( A167  and  (not A169) );
 a287a <=( (not a285a)  and  (not a286a) );
 a288a <=( A166  and  (not a287a) );
 a289a <=( (not A170)  and  (not a51a) );
 a290a <=( A169  and  (not a289a) );
 a291a <=( (not A169)  and  (not A170) );
 a292a <=( (not a290a)  and  (not a291a) );
 a293a <=( (not a288a)  and  a292a );
 a294a <=( (not A168)  and  (not a293a) );
 a295a <=( a83a  and  (not a264a) );
 a296a <=( (not a294a)  and  (not a295a) );
 a297a <=( (not a284a)  and  (not a296a) );
 a298a <=( A234  and  a116a );
 a299a <=( (not a95a)  and  a298a );
 a300a <=( (not a117a)  and  (not a299a) );
 a301a <=( A267  and  A265 );
 a302a <=( (not a108a)  and  a301a );
 a303a <=( (not A266)  and  (not a302a) );
 a304a <=( (not a122a)  and  (not a303a) );
 a305a <=( A300  and  A298 );
 a306a <=( (not a99a)  and  a305a );
 a307a <=( (not A299)  and  (not a306a) );
 a308a <=( (not a130a)  and  (not a307a) );
 a309a <=( (not a304a)  and  (not a308a) );
 a310a <=( (not a300a)  and  a309a );
 a311a <=( (not a263a)  and  (not a310a) );
 a312a <=( (not a280a)  and  a311a );
 A109 <=( (not a297a)  and  a312a );
 a314a <=( (not a55a)  and  (not a143a) );
 a315a <=( (not a254a)  and  a314a );
 a316a <=( (not a278a)  and  a315a );
 a317a <=( (not a309a)  and  a316a );
 a318a <=( (not a276a)  and  (not a317a) );
 A108 <=( (not a297a)  and  (not a318a) );
 a320a <=( (not a96a)  and  (not a257a) );
 a321a <=( (not a296a)  and  (not a320a) );
 a322a <=( a300a  and  (not a321a) );
 a323a <=( (not a279a)  and  (not a322a) );
 a324a <=( (not a284a)  and  (not a320a) );
 a325a <=( a300a  and  (not a324a) );
 a326a <=( (not a276a)  and  (not a325a) );
 a327a <=( (not a105a)  and  (not a259a) );
 a328a <=( (not a326a)  and  a327a );
 a329a <=( (not a323a)  and  a328a );
 a330a <=( (not a308a)  and  (not a327a) );
 a331a <=( (not a276a)  and  a330a );
 a332a <=( (not a304a)  and  (not a320a) );
 a333a <=( (not a296a)  and  a332a );
 a334a <=( a300a  and  (not a331a) );
 a335a <=( (not a333a)  and  a334a );
 a336a <=( (not a279a)  and  (not a335a) );
 a337a <=( (not a284a)  and  (not a304a) );
 a338a <=( (not a320a)  and  a337a );
 a339a <=( a300a  and  (not a338a) );
 a340a <=( (not a276a)  and  (not a339a) );
 a341a <=( (not a284a)  and  (not a308a) );
 a342a <=( (not a327a)  and  a341a );
 a343a <=( (not a296a)  and  a342a );
 a344a <=( (not a340a)  and  (not a343a) );
 a345a <=( (not a336a)  and  a344a );
 a346a <=( (not a105a)  and  (not a130a) );
 a347a <=( (not a307a)  and  a346a );
 a348a <=( (not a259a)  and  a347a );
 a349a <=( (not a255a)  and  (not a348a) );
 a350a <=( (not a300a)  and  a332a );
 a351a <=( (not a349a)  and  (not a350a) );
 a352a <=( (not a280a)  and  a351a );
 A105 <=( (not a297a)  and  a352a );
 a354a <=( A236  and  (not a142a) );
 a355a <=( (not A234)  and  (not a354a) );
 a356a <=( (not a143a)  and  (not a355a) );
 a357a <=( A302  and  (not a98a) );
 a358a <=( A300  and  (not a131a) );
 a359a <=( A269  and  (not a107a) );
 a360a <=( A267  and  (not a123a) );
 a361a <=( (not A301)  and  (not A268) );
 a362a <=( (not a360a)  and  a361a );
 a363a <=( (not a358a)  and  a362a );
 a364a <=( (not a357a)  and  (not a359a) );
 a365a <=( a363a  and  a364a );
 a366a <=( (not A235)  and  (not a356a) );
 a367a <=( (not a365a)  and  a366a );
 a368a <=( A170  and  (not a82a) );
 a369a <=( (not A168)  and  (not a368a) );
 a370a <=( (not a83a)  and  (not a369a) );
 a371a <=( A203  and  (not a68a) );
 a372a <=( (not A201)  and  (not a371a) );
 a373a <=( (not a69a)  and  (not a372a) );
 a374a <=( (not A202)  and  (not A169) );
 a375a <=( (not a373a)  and  a374a );
 a376a <=( (not a370a)  and  a375a );
 a377a <=( (not A167)  and  A170 );
 a378a <=( (not A168)  and  (not a377a) );
 a379a <=( A166  and  (not a378a) );
 a380a <=( (not A166)  and  A170 );
 a381a <=( (not A168)  and  (not a380a) );
 a382a <=( A167  and  (not a381a) );
 a383a <=( (not A169)  and  (not a382a) );
 a384a <=( (not a379a)  and  a383a );
 a385a <=( A203  and  (not a56a) );
 a386a <=( A201  and  (not a69a) );
 a387a <=( (not A202)  and  (not a386a) );
 a388a <=( (not a385a)  and  a387a );
 a389a <=( (not a384a)  and  (not a388a) );
 a390a <=( A269  and  (not a122a) );
 a391a <=( (not A267)  and  (not a390a) );
 a392a <=( (not a123a)  and  (not a391a) );
 a393a <=( A302  and  (not a130a) );
 a394a <=( (not A300)  and  (not a393a) );
 a395a <=( (not a131a)  and  (not a394a) );
 a396a <=( A236  and  (not a118a) );
 a397a <=( A234  and  (not a143a) );
 a398a <=( (not A235)  and  (not a397a) );
 a399a <=( (not a396a)  and  a398a );
 a400a <=( a361a  and  (not a399a) );
 a401a <=( (not a392a)  and  (not a395a) );
 a402a <=( a400a  and  a401a );
 a403a <=( (not a389a)  and  (not a402a) );
 a404a <=( (not a367a)  and  (not a376a) );
 A76 <=( a403a  and  a404a );
 a406a <=( a361a  and  (not a395a) );
 a407a <=( (not a392a)  and  a406a );
 a408a <=( (not a366a)  and  a388a );
 a409a <=( (not a407a)  and  a408a );
 a410a <=( (not a384a)  and  (not a409a) );
 A75 <=( (not a376a)  and  (not a410a) );
 a412a <=( (not A301)  and  (not a358a) );
 a413a <=( (not a357a)  and  a412a );
 a414a <=( (not A169)  and  (not a413a) );
 a415a <=( (not a370a)  and  a414a );
 a416a <=( a399a  and  (not a415a) );
 a417a <=( (not a388a)  and  (not a416a) );
 a418a <=( (not A202)  and  (not a413a) );
 a419a <=( (not a373a)  and  a418a );
 a420a <=( a399a  and  (not a419a) );
 a421a <=( (not a384a)  and  (not a420a) );
 a422a <=( (not A268)  and  (not a360a) );
 a423a <=( (not a359a)  and  a422a );
 a424a <=( (not a421a)  and  a423a );
 a425a <=( (not a417a)  and  a424a );
 a426a <=( (not a392a)  and  (not a413a) );
 a427a <=( (not A268)  and  (not A169) );
 a428a <=( (not a370a)  and  a427a );
 a429a <=( a426a  and  a428a );
 a430a <=( (not A301)  and  (not a423a) );
 a431a <=( (not a395a)  and  a430a );
 a432a <=( (not a384a)  and  a431a );
 a433a <=( a399a  and  (not a429a) );
 a434a <=( (not a432a)  and  a433a );
 a435a <=( (not a388a)  and  (not a434a) );
 a436a <=( (not A268)  and  (not A202) );
 a437a <=( (not a373a)  and  a436a );
 a438a <=( a426a  and  a437a );
 a439a <=( a399a  and  (not a438a) );
 a440a <=( (not a384a)  and  (not a439a) );
 a441a <=( (not A301)  and  a374a );
 a442a <=( (not a423a)  and  a441a );
 a443a <=( (not a373a)  and  (not a395a) );
 a444a <=( (not a370a)  and  a443a );
 a445a <=( a442a  and  a444a );
 a446a <=( (not a440a)  and  (not a445a) );
 a447a <=( (not a435a)  and  a446a );
 a448a <=( (not A301)  and  (not a395a) );
 a449a <=( a423a  and  (not a448a) );
 a450a <=( a366a  and  (not a449a) );
 a451a <=( (not A268)  and  (not a413a) );
 a452a <=( (not a392a)  and  (not a399a) );
 a453a <=( a451a  and  a452a );
 a454a <=( (not a389a)  and  (not a453a) );
 a455a <=( (not a376a)  and  a454a );
 A72 <=( (not a450a)  and  a455a );
 a457a <=( (not A203)  and  A202 );
 a458a <=( (not a70a)  and  a457a );
 a459a <=( (not A202)  and  a385a );
 a460a <=( (not a386a)  and  (not a458a) );
 a461a <=( (not a459a)  and  a460a );
 a462a <=( A168  and  (not a291a) );
 a463a <=( a52a  and  a462a );
 a464a <=( (not a51a)  and  (not a463a) );
 a465a <=( (not a461a)  and  (not a464a) );
 a466a <=( A166  and  a462a );
 a467a <=( (not A167)  and  (not a466a) );
 a468a <=( (not a82a)  and  (not a467a) );
 a469a <=( A203  and  (not A202) );
 a470a <=( (not a56a)  and  (not a469a) );
 a471a <=( a68a  and  (not a457a) );
 a472a <=( (not a470a)  and  (not a471a) );
 a473a <=( (not a468a)  and  (not a472a) );
 a474a <=( (not A201)  and  a473a );
 a475a <=( a69a  and  (not a457a) );
 a476a <=( (not a468a)  and  a475a );
 a477a <=( A236  and  (not A235) );
 a478a <=( (not A302)  and  A301 );
 a479a <=( (not a132a)  and  a478a );
 a480a <=( (not A301)  and  a357a );
 a481a <=( (not A269)  and  A268 );
 a482a <=( (not a124a)  and  a481a );
 a483a <=( (not A268)  and  a359a );
 a484a <=( (not a360a)  and  (not a482a) );
 a485a <=( (not a483a)  and  a484a );
 a486a <=( (not a358a)  and  (not a479a) );
 a487a <=( (not a480a)  and  a486a );
 a488a <=( a485a  and  a487a );
 a489a <=( (not A234)  and  (not a477a) );
 a490a <=( (not a488a)  and  a489a );
 a491a <=( A269  and  (not A268) );
 a492a <=( A302  and  (not A301) );
 a493a <=( (not a98a)  and  (not a492a) );
 a494a <=( a130a  and  (not a478a) );
 a495a <=( (not a493a)  and  (not a494a) );
 a496a <=( (not a107a)  and  (not a491a) );
 a497a <=( (not a495a)  and  a496a );
 a498a <=( a122a  and  (not a481a) );
 a499a <=( (not a495a)  and  a498a );
 a500a <=( (not a497a)  and  (not a499a) );
 a501a <=( (not A300)  and  (not a500a) );
 a502a <=( (not a496a)  and  (not a498a) );
 a503a <=( a131a  and  (not a478a) );
 a504a <=( (not a502a)  and  a503a );
 a505a <=( (not a501a)  and  (not a504a) );
 a506a <=( (not A267)  and  (not a505a) );
 a507a <=( (not A300)  and  (not a495a) );
 a508a <=( (not a503a)  and  (not a507a) );
 a509a <=( a123a  and  (not a481a) );
 a510a <=( (not a508a)  and  a509a );
 a511a <=( (not a506a)  and  (not a510a) );
 a512a <=( a477a  and  (not a511a) );
 a513a <=( (not a490a)  and  (not a512a) );
 a514a <=( (not a118a)  and  (not a513a) );
 a515a <=( (not A234)  and  a142a );
 a516a <=( (not a143a)  and  (not a515a) );
 a517a <=( (not A236)  and  A235 );
 a518a <=( (not a516a)  and  (not a517a) );
 a519a <=( (not a488a)  and  a518a );
 a520a <=( (not a144a)  and  a517a );
 a521a <=( (not a397a)  and  (not a520a) );
 a522a <=( (not A300)  and  (not a521a) );
 a523a <=( (not a500a)  and  a522a );
 a524a <=( (not a502a)  and  (not a521a) );
 a525a <=( a503a  and  a524a );
 a526a <=( (not a523a)  and  (not a525a) );
 a527a <=( (not A267)  and  (not a526a) );
 a528a <=( (not a495a)  and  a522a );
 a529a <=( a503a  and  (not a521a) );
 a530a <=( (not a528a)  and  (not a529a) );
 a531a <=( a509a  and  (not a530a) );
 a532a <=( (not a465a)  and  (not a476a) );
 a533a <=( (not a519a)  and  a532a );
 a534a <=( (not a474a)  and  a533a );
 a535a <=( (not a531a)  and  a534a );
 a536a <=( (not a527a)  and  a535a );
 A43 <=( (not a514a)  and  a536a );
 a538a <=( (not a118a)  and  (not a477a) );
 a539a <=( a142a  and  (not a517a) );
 a540a <=( (not a538a)  and  (not a539a) );
 a541a <=( (not A234)  and  (not a540a) );
 a542a <=( (not a464a)  and  a541a );
 a543a <=( a143a  and  (not a517a) );
 a544a <=( (not a386a)  and  (not a543a) );
 a545a <=( (not a458a)  and  a544a );
 a546a <=( (not a459a)  and  a545a );
 a547a <=( a511a  and  a546a );
 a548a <=( (not a464a)  and  (not a547a) );
 a549a <=( (not a476a)  and  (not a542a) );
 a550a <=( (not a474a)  and  a549a );
 A42 <=( (not a548a)  and  a550a );
 a552a <=( (not A235)  and  a396a );
 a553a <=( a521a  and  (not a552a) );
 a554a <=( a460a  and  a464a );
 a555a <=( (not a459a)  and  a554a );
 a556a <=( (not a553a)  and  (not a555a) );
 a557a <=( (not a468a)  and  (not a487a) );
 a558a <=( (not a461a)  and  a557a );
 a559a <=( (not a464a)  and  (not a472a) );
 a560a <=( (not a487a)  and  a559a );
 a561a <=( (not A201)  and  a560a );
 a562a <=( (not a464a)  and  (not a487a) );
 a563a <=( a475a  and  a562a );
 a564a <=( a485a  and  (not a563a) );
 a565a <=( (not a558a)  and  (not a561a) );
 a566a <=( (not a556a)  and  a565a );
 a567a <=( a564a  and  a566a );
 a568a <=( (not a464a)  and  a507a );
 a569a <=( (not a464a)  and  a503a );
 a570a <=( (not a568a)  and  (not a569a) );
 a571a <=( (not a485a)  and  (not a570a) );
 a572a <=( (not A267)  and  (not a502a) );
 a573a <=( (not a468a)  and  a572a );
 a574a <=( (not a487a)  and  a573a );
 a575a <=( a509a  and  a557a );
 a576a <=( (not a574a)  and  (not a575a) );
 a577a <=( (not a571a)  and  a576a );
 a578a <=( (not a461a)  and  (not a577a) );
 a579a <=( (not A300)  and  a491a );
 a580a <=( (not a492a)  and  a579a );
 a581a <=( a473a  and  a580a );
 a582a <=( A302  and  (not A267) );
 a583a <=( (not A301)  and  a582a );
 a584a <=( (not a491a)  and  a583a );
 a585a <=( a559a  and  a584a );
 a586a <=( (not a581a)  and  (not a585a) );
 a587a <=( (not a98a)  and  (not a586a) );
 a588a <=( (not A300)  and  a130a );
 a589a <=( (not a131a)  and  (not a588a) );
 a590a <=( (not a478a)  and  a491a );
 a591a <=( (not a589a)  and  a590a );
 a592a <=( a473a  and  a591a );
 a593a <=( (not A267)  and  (not a491a) );
 a594a <=( (not a486a)  and  a593a );
 a595a <=( a559a  and  a594a );
 a596a <=( (not a592a)  and  (not a595a) );
 a597a <=( (not a587a)  and  a596a );
 a598a <=( (not a107a)  and  (not a597a) );
 a599a <=( (not A267)  and  a122a );
 a600a <=( (not a123a)  and  (not a599a) );
 a601a <=( (not a481a)  and  (not a600a) );
 a602a <=( a560a  and  a601a );
 a603a <=( a470a  and  (not a495a) );
 a604a <=( a471a  and  (not a495a) );
 a605a <=( (not a603a)  and  (not a604a) );
 a606a <=( (not A300)  and  (not a484a) );
 a607a <=( (not a468a)  and  a606a );
 a608a <=( (not a605a)  and  a607a );
 a609a <=( (not a484a)  and  a503a );
 a610a <=( (not a472a)  and  a609a );
 a611a <=( (not a468a)  and  a610a );
 a612a <=( (not a608a)  and  (not a611a) );
 a613a <=( (not a602a)  and  a612a );
 a614a <=( (not a598a)  and  a613a );
 a615a <=( (not A201)  and  (not a614a) );
 a616a <=( (not a468a)  and  a580a );
 a617a <=( (not a464a)  and  a584a );
 a618a <=( (not a616a)  and  (not a617a) );
 a619a <=( (not a98a)  and  (not a618a) );
 a620a <=( (not a468a)  and  a591a );
 a621a <=( (not a464a)  and  a594a );
 a622a <=( (not a620a)  and  (not a621a) );
 a623a <=( (not a619a)  and  a622a );
 a624a <=( (not a107a)  and  (not a623a) );
 a625a <=( a562a  and  a601a );
 a626a <=( (not a495a)  and  a606a );
 a627a <=( (not a468a)  and  a626a );
 a628a <=( (not a468a)  and  a609a );
 a629a <=( (not a627a)  and  (not a628a) );
 a630a <=( (not a625a)  and  a629a );
 a631a <=( (not a624a)  and  a630a );
 a632a <=( a475a  and  (not a631a) );
 a633a <=( (not a556a)  and  (not a578a) );
 a634a <=( (not a632a)  and  a633a );
 a635a <=( (not a615a)  and  a634a );
 a636a <=( a485a  and  (not a503a) );
 a637a <=( (not a507a)  and  a636a );
 a638a <=( a489a  and  (not a637a) );
 a639a <=( (not a487a)  and  a572a );
 a640a <=( (not a487a)  and  a509a );
 a641a <=( (not a639a)  and  (not a640a) );
 a642a <=( a477a  and  (not a641a) );
 a643a <=( (not a638a)  and  (not a642a) );
 a644a <=( (not a118a)  and  (not a643a) );
 a645a <=( a518a  and  (not a637a) );
 a646a <=( (not A267)  and  (not a487a) );
 a647a <=( a524a  and  a646a );
 a648a <=( a509a  and  (not a521a) );
 a649a <=( (not a487a)  and  a648a );
 a650a <=( (not a476a)  and  (not a649a) );
 a651a <=( (not a465a)  and  a650a );
 a652a <=( (not a474a)  and  (not a647a) );
 a653a <=( a651a  and  a652a );
 a654a <=( (not a645a)  and  a653a );
 A39 <=( (not a644a)  and  a654a );
 a656a <=( A300  and  (not a492a) );
 a657a <=( A302  and  (not A300) );
 a658a <=( (not A301)  and  a657a );
 a659a <=( (not a656a)  and  (not a658a) );
 a660a <=( (not a98a)  and  (not a107a) );
 a661a <=( (not a659a)  and  a660a );
 a662a <=( A267  and  a661a );
 a663a <=( (not A300)  and  (not a492a) );
 a664a <=( A302  and  A300 );
 a665a <=( (not A301)  and  a664a );
 a666a <=( a132a  and  (not a665a) );
 a667a <=( (not a663a)  and  a666a );
 a668a <=( (not A267)  and  (not a667a) );
 a669a <=( (not a662a)  and  (not a668a) );
 a670a <=( (not a491a)  and  (not a669a) );
 a671a <=( (not A267)  and  (not a107a) );
 a672a <=( (not a98a)  and  a671a );
 a673a <=( A300  and  a672a );
 a674a <=( (not A300)  and  A267 );
 a675a <=( (not a673a)  and  (not a674a) );
 a676a <=( a491a  and  (not a675a) );
 a677a <=( (not A300)  and  (not a124a) );
 a678a <=( (not a676a)  and  (not a677a) );
 a679a <=( (not a492a)  and  (not a678a) );
 a680a <=( A269  and  A267 );
 a681a <=( (not A268)  and  a680a );
 a682a <=( a124a  and  (not a681a) );
 a683a <=( (not a666a)  and  (not a682a) );
 a684a <=( a491a  and  a658a );
 a685a <=( a672a  and  a684a );
 a686a <=( A201  and  (not a469a) );
 a687a <=( A203  and  (not A201) );
 a688a <=( (not A202)  and  a687a );
 a689a <=( (not a686a)  and  (not a688a) );
 a690a <=( (not a56a)  and  (not a689a) );
 a691a <=( (not A168)  and  (not a291a) );
 a692a <=( A168  and  a291a );
 a693a <=( a84a  and  (not a692a) );
 a694a <=( (not a691a)  and  a693a );
 a695a <=( (not a690a)  and  a694a );
 a696a <=( (not A234)  and  (not a695a) );
 a697a <=( (not A168)  and  a291a );
 a698a <=( (not a462a)  and  (not a697a) );
 a699a <=( (not A201)  and  (not a469a) );
 a700a <=( A203  and  A201 );
 a701a <=( (not A202)  and  a700a );
 a702a <=( a70a  and  (not a701a) );
 a703a <=( (not a699a)  and  a702a );
 a704a <=( A234  and  (not a118a) );
 a705a <=( (not a53a)  and  a704a );
 a706a <=( (not a698a)  and  a705a );
 a707a <=( (not a703a)  and  a706a );
 a708a <=( (not a696a)  and  (not a707a) );
 a709a <=( (not a477a)  and  (not a708a) );
 a710a <=( A236  and  A234 );
 a711a <=( (not A235)  and  a710a );
 a712a <=( a144a  and  (not a711a) );
 a713a <=( (not a56a)  and  (not a712a) );
 a714a <=( (not a689a)  and  a713a );
 a715a <=( (not A168)  and  (not a712a) );
 a716a <=( (not a53a)  and  (not a118a) );
 a717a <=( (not a703a)  and  a716a );
 a718a <=( (not A234)  and  A168 );
 a719a <=( a477a  and  a718a );
 a720a <=( a717a  and  a719a );
 a721a <=( (not a715a)  and  (not a720a) );
 a722a <=( (not a291a)  and  (not a721a) );
 a723a <=( (not a693a)  and  (not a712a) );
 a724a <=( (not A234)  and  (not A168) );
 a725a <=( a477a  and  a724a );
 a726a <=( a291a  and  a725a );
 a727a <=( a717a  and  a726a );
 a728a <=( (not a683a)  and  (not a723a) );
 a729a <=( (not a714a)  and  a728a );
 a730a <=( (not a685a)  and  a729a );
 a731a <=( (not a727a)  and  a730a );
 a732a <=( (not a670a)  and  a731a );
 a733a <=( (not a709a)  and  (not a722a) );
 a734a <=( a732a  and  a733a );
 A6 <=( (not a679a)  and  a734a );
 a736a <=( (not a53a)  and  (not a698a) );
 a737a <=( a703a  and  (not a736a) );
 a738a <=( (not A267)  and  (not a737a) );
 a739a <=( (not a489a)  and  a712a );
 a740a <=( (not a694a)  and  (not a739a) );
 a741a <=( A267  and  (not a107a) );
 a742a <=( a740a  and  a741a );
 a743a <=( (not a738a)  and  (not a742a) );
 a744a <=( (not A300)  and  (not a743a) );
 a745a <=( (not a53a)  and  (not a107a) );
 a746a <=( A267  and  A168 );
 a747a <=( a745a  and  a746a );
 a748a <=( (not a188a)  and  (not a747a) );
 a749a <=( (not a291a)  and  (not a739a) );
 a750a <=( (not a748a)  and  a749a );
 a751a <=( A267  and  (not A168) );
 a752a <=( a745a  and  a751a );
 a753a <=( (not A267)  and  A168 );
 a754a <=( (not a752a)  and  (not a753a) );
 a755a <=( a291a  and  (not a754a) );
 a756a <=( (not A267)  and  (not a84a) );
 a757a <=( (not a755a)  and  (not a756a) );
 a758a <=( (not a739a)  and  (not a757a) );
 a759a <=( (not a750a)  and  (not a758a) );
 a760a <=( (not a98a)  and  (not a759a) );
 a761a <=( A300  and  a760a );
 a762a <=( (not a744a)  and  (not a761a) );
 a763a <=( (not a492a)  and  (not a762a) );
 a764a <=( (not a666a)  and  (not a743a) );
 a765a <=( a658a  and  a760a );
 a766a <=( (not a764a)  and  (not a765a) );
 a767a <=( (not a763a)  and  a766a );
 a768a <=( (not a491a)  and  (not a767a) );
 a769a <=( (not A300)  and  (not a737a) );
 a770a <=( (not a98a)  and  a740a );
 a771a <=( A300  and  a770a );
 a772a <=( (not a769a)  and  (not a771a) );
 a773a <=( (not a492a)  and  (not a772a) );
 a774a <=( (not a666a)  and  (not a737a) );
 a775a <=( a658a  and  a770a );
 a776a <=( (not a774a)  and  (not a775a) );
 a777a <=( (not a773a)  and  a776a );
 a778a <=( (not a682a)  and  (not a777a) );
 a779a <=( a690a  and  (not a739a) );
 a780a <=( A269  and  (not A267) );
 a781a <=( (not A268)  and  a780a );
 a782a <=( (not a98a)  and  a781a );
 a783a <=( (not a107a)  and  a782a );
 a784a <=( (not a659a)  and  a783a );
 a785a <=( (not a739a)  and  a784a );
 a786a <=( (not a779a)  and  (not a785a) );
 a787a <=( a63a  and  (not a786a) );
 a788a <=( (not a107a)  and  a781a );
 a789a <=( (not a667a)  and  a788a );
 a790a <=( a703a  and  (not a789a) );
 a791a <=( (not A168)  and  (not a739a) );
 a792a <=( (not a790a)  and  a791a );
 a793a <=( (not a787a)  and  (not a792a) );
 a794a <=( (not a291a)  and  (not a793a) );
 a795a <=( a661a  and  a781a );
 a796a <=( (not a690a)  and  (not a795a) );
 a797a <=( (not A168)  and  (not a53a) );
 a798a <=( (not a796a)  and  a797a );
 a799a <=( A168  and  (not a790a) );
 a800a <=( (not a798a)  and  (not a799a) );
 a801a <=( a291a  and  (not a800a) );
 a802a <=( (not a84a)  and  (not a790a) );
 a803a <=( (not a801a)  and  (not a802a) );
 a804a <=( (not a739a)  and  (not a803a) );
 a805a <=( (not a794a)  and  (not a804a) );
 a806a <=( (not a778a)  and  a805a );
 A7 <=( (not a768a)  and  a806a );
 a808a <=( A234  and  (not a477a) );
 a809a <=( A236  and  (not A234) );
 a810a <=( (not A235)  and  a809a );
 a811a <=( (not a808a)  and  (not a810a) );
 a812a <=( (not a98a)  and  (not a811a) );
 a813a <=( (not a659a)  and  a812a );
 a814a <=( A267  and  (not a491a) );
 a815a <=( (not a781a)  and  (not a814a) );
 a816a <=( (not a107a)  and  (not a815a) );
 a817a <=( (not a811a)  and  a816a );
 a818a <=( (not a813a)  and  (not a817a) );
 a819a <=( (not a118a)  and  (not a818a) );
 a820a <=( (not a593a)  and  a682a );
 a821a <=( (not a98a)  and  (not a659a) );
 a822a <=( (not a820a)  and  a821a );
 a823a <=( (not a667a)  and  a816a );
 a824a <=( (not a822a)  and  (not a823a) );
 a825a <=( a736a  and  (not a824a) );
 a826a <=( (not a690a)  and  (not a825a) );
 a827a <=( (not a819a)  and  a826a );
 a828a <=( (not a694a)  and  (not a703a) );
 a829a <=( (not a489a)  and  (not a663a) );
 a830a <=( a712a  and  a829a );
 a831a <=( a666a  and  a830a );
 a832a <=( (not a828a)  and  a831a );
 a833a <=( (not A267)  and  (not a832a) );
 a834a <=( (not a662a)  and  (not a833a) );
 a835a <=( (not a491a)  and  (not a834a) );
 a836a <=( (not a682a)  and  (not a832a) );
 a837a <=( (not a795a)  and  (not a836a) );
 A9 <=( (not a835a)  and  a837a );
 a839a <=( (not a690a)  and  (not a736a) );
 a840a <=( (not A234)  and  (not a839a) );
 a841a <=( (not a118a)  and  a828a );
 a842a <=( A234  and  a841a );
 a843a <=( (not a840a)  and  (not a842a) );
 a844a <=( (not a477a)  and  (not a843a) );
 a845a <=( (not a53a)  and  (not a712a) );
 a846a <=( (not a698a)  and  a845a );
 a847a <=( a810a  and  a841a );
 a848a <=( (not a683a)  and  (not a846a) );
 a849a <=( (not a685a)  and  (not a714a) );
 a850a <=( a848a  and  a849a );
 a851a <=( (not a847a)  and  a850a );
 a852a <=( (not a670a)  and  a851a );
 a853a <=( (not a844a)  and  a852a );
 A10 <=( (not a679a)  and  a853a );
 A140 <=( (not a187a) );
 A139 <=( (not a221a) );
 A107 <=( (not a329a) );
 A106 <=( (not a345a) );
 A74 <=( (not a425a) );
 A73 <=( (not a447a) );
 A41 <=( (not a567a) );
 A40 <=( (not a635a) );
 A8 <=( (not a827a) );


end testing_behav;
